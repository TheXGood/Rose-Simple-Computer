module controlunit(clk);

	input wire clk;
	
	
	

end