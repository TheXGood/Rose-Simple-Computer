//Interrupt Controller

module InterruptController(clk,IntNo,Except,);
	
	
endmodule